-- Hassanal Harriz Bin Ahmed Hakimmy Fuad
-- U2102848

library ieee;
use ieee.std_logic_1164.all;

use work.components.all;

entity sort is
	generic ( N : integer := 8 );
	
	port ( 	Clock, ResetN  	: IN     STD_LOGIC;
			S, WrInit, Rd 	: IN     STD_LOGIC;
			DataIn			: IN 	 STD_LOGIC_VECTOR (N-1 downto 0);
			RAdd			: IN 	 integer range 0 to N-1;
			DataOut			: BUFFER STD_LOGIC_VECTOR (N-1 downto 0);
			Done			: BUFFER STD_LOGIC
		);

end sort;

architecture dataflow of sort is

-- datapath data buses
	type RegArray is ARRAY (7 downto 0) of STD_LOGIC_VECTOR (N-1 downto 0);
	signal R 		: RegArray;
	signal RData	: STD_LOGIC_VECTOR (N-1 downto 0);
	signal ABData	: STD_LOGIC_VECTOR (N-1 downto 0);
	signal A, B 	: STD_LOGIC_VECTOR (N-1 downto 0);
	signal ABMux	: STD_LOGIC_VECTOR (N-1 downto 0);
	
-- datapath control signals
	signal Rin			: STD_LOGIC_VECTOR (7 downto 0);
	signal IMux			: integer range 0 to 7;
	signal Ain, Bin		: STD_LOGIC;
	signal Aout, Bout	: STD_LOGIC;
	signal BItA			: STD_LOGIC;

-- control unit Part 1
	signal Zero			: integer range 7 downto 0;
	signal Ci, Cj		: integer range 0 to 7;
	signal CMux			: integer range 0 to 7;
	
	signal LI, LJ		: STD_LOGIC;
	signal EI, EJ		: STD_LOGIC;
	
	signal zi, zj		: STD_LOGIC;
	signal Csel			: STD_LOGIC;
	signal Int			: STD_LOGIC;
	signal Wr			: STD_LOGIC;

-- control unit Part 2
	type State_type is ( S1, S2, S3, S4, S5, S6, S7, S8, S9 );
	signal y : State_type;
	

begin 
	RData <= ABMux when WrInit = '0' else DataIn;
	
	GenReg: for i in 0 to 7 generate
		Reg: registEn generic map ( N => N )
		port map (	D		=> RData,
					ResetN	=> ResetN,
					E 		=> Rin(i),
					Clock 	=> Clock,
					Q		=> R(i)
				);
	end generate;
	
	with IMux select
		ABData <= 	R(0) when 0,
					R(1) when 1,
					R(2) when 2,
					R(3) when 3,
					R(4) when 4,
					R(5) when 5,
					R(6) when 6,
					R(7) when others;
					
	RegA: registEn generic map ( N => N )
		port map (	D		=> ABData,
					ResetN	=> ResetN,
					E 		=> Ain,
					Clock 	=> Clock,
					Q		=> A
				);
	
	RegB: registEn generic map ( N => N )
		port map (	D		=> ABData,
					ResetN	=> ResetN,
					E 		=> Bin,
					Clock 	=> Clock,
					Q		=> B
				);
	
	BItA <= '1' when B < A else '0';
	ABMux <= A when Bout = '0' else B;
	DataOut <= (others => 'Z') when Rd = '0' else ABData;
	
	Zero <= 0;
	OuterLoop : upcount generic map ( modulus => 8 )
		port map (	ResetN	=> ResetN,
					Clock	=> Clock,
					E		=> EI,
					L		=> LI,
					R		=> Zero,
					Q		=> Ci
				);
	
	InnerLoop : upcount generic map ( modulus => 8 )
		port map (	ResetN	=> ResetN,
					Clock	=> Clock,
					E		=> EJ,
					L		=> LJ,
					R		=> Ci,
					Q		=> Cj
				);
	
	CMux <= Ci when Csel = '0' else Cj;
	IMux <= CMux when Int = '1' else RAdd;
	
	
	RinDec: process (WrInit, Wr, IMux)
	begin
		if (WrInit or Wr) = '1' then
			case IMux is
				when 0		=> Rin <= "00000001";
				when 1		=> Rin <= "00000010";
				when 2		=> Rin <= "00000100";
				when 3		=> Rin <= "00001000";
				when 4		=> Rin <= "00010000";
				when 5		=> Rin <= "00100000";
				when 6		=> Rin <= "01000000";
				when others	=> Rin <= "10000000";
			end case;
		else Rin <= "00000000";
		end if;
	end process;
	
	zi <= '1' when Ci = 6 else '0';
	zj <= '1' when Cj = 7 else '0';
	

	FSM_transitions: process (ResetN, Clock)
		begin
			if ResetN = '0' then
				y <= S1;
			elsif (Clock'EVENT and Clock = '1' ) then 
				case y is
					when S1		=> 	if S = '0' then y <= S1; else y <= S2; end if;
									
					when S2		=> 	y <= S3;
					
					when S3		=> 	y <= S4;
					
					when S4		=> 	y <= S5;
					
					when S5		=> 	if BItA = '1' then y <= S6; else y <= S8; end if;
					
					when S6		=> 	y <= S7;
					
					when S7		=> 	y <= S8;
					
					when S8		=>	if zj = '0' then y <= S4; elsif zi = '0' then y <= S2; else y <= S9; end if;
					
					when others	=> 	if S = '1' then y <= S9; else y <= S1; end if;
				end case;
			end if;
	end process;
	
-- define the outputs generated by the FSM
	Int <= '0'	when y = S1		else '1';
	Done <= '1'	when y = S9		else '0';
	
	FSM_outputs: process (y, zi, zj)
	begin
		LI 		<= '0';
		LJ 		<= '0';
		EI 		<= '0';
		EJ 		<= '0';
		Csel 	<= '0';
		Wr 		<= '0';
		Ain 	<= '0';
		Bin 	<= '0';
		Aout 	<= '0';
		Bout 	<= '0';
		case y is
			when S1		=> LI <= '1'; EI <= '1';
			when S2		=> Ain <= '1'; LJ <= '1'; EJ <= '1';
			when S3		=> EJ <= '1';
			when S4		=> Bin <= '1'; Csel <= '1';
			when S5		=> -- no outputs asserted in this state
			when S6		=> Csel <= '1'; Wr <= '1'; Aout <= '1';
			when S7		=> Wr <= '1'; Bout <= '1';
			when S8		=>	Ain <= '1';
							if zj = '0' then 
								EJ <= '1';
							else
								EJ <= '0';
								if zi = '0' then 
									EI <= '1';
								else
									EI <= '0';
								end if;
							end if;
			when others	=> -- Done is assigned 1 by conditional signal assignment
		end case;
	end process;
	
end dataflow;