-- Hassanal Harriz Bin Ahmed Hakimmy Fuad
-- U2102848

library ieee;
use ieee.std_logic_1164.all;

entity DFF is
	port (	din		: in  std_logic;
			clk		: in  std_logic;
			rst		: in  std_logic;
			dout	: out std_logic
		);
end DFF;

architecture behavioral of DFF is 
begin
	process (rst, clk, din)
	begin
		if (rst ='1') then 
			dout <= '0';
		elsif (rising_edge(clk)) then
			dout <= din;
		end if;
	end process;
end architecture;